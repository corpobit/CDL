---logs:[t:timestamp:time|n:temp|n:humidity:1623456789,23.5,45.2,1623456790,24.1,44.8]---
