---company:(
  name|departments:
  "MegaCorp",
  [name|employees:
    Engineering,[name|role:
      Employee1,Engineer,
      Employee2,Engineer,
      Employee3,Engineer,
      Employee4,Engineer,
      Employee5,Engineer,
      Employee6,Engineer,
      Employee7,Engineer,
      Employee8,Engineer,
      Employee9,Engineer,
      Employee10,Engineer,
      Employee11,Engineer,
      Employee12,Engineer,
      Employee13,Engineer,
      Employee14,Engineer,
      Employee15,Engineer,
      Employee16,Engineer,
      Employee17,Engineer,
      Employee18,Engineer,
      Employee19,Engineer,
      Employee20,Engineer,
      Employee21,Engineer,
      Employee22,Engineer,
      Employee23,Engineer,
      Employee24,Engineer,
      Employee25,Engineer,
      Employee26,Engineer,
      Employee27,Engineer,
      Employee28,Engineer,
      Employee29,Engineer,
      Employee30,Engineer,
      Employee31,Engineer,
      Employee32,Engineer,
      Employee33,Engineer,
      Employee34,Engineer,
      Employee35,Engineer,
      Employee36,Engineer,
      Employee37,Engineer,
      Employee38,Engineer,
      Employee39,Engineer,
      Employee40,Engineer,
      Employee41,Engineer,
      Employee42,Engineer,
      Employee43,Engineer,
      Employee44,Engineer,
      Employee45,Engineer,
      Employee46,Engineer,
      Employee47,Engineer,
      Employee48,Engineer,
      Employee49,Engineer,
      Employee50,Engineer,
      Employee51,Engineer,
      Employee52,Engineer,
      Employee53,Engineer,
      Employee54,Engineer,
      Employee55,Engineer,
      Employee56,Engineer,
      Employee57,Engineer,
      Employee58,Engineer,
      Employee59,Engineer,
      Employee60,Engineer,
      Employee61,Engineer,
      Employee62,Engineer,
      Employee63,Engineer,
      Employee64,Engineer,
      Employee65,Engineer,
      Employee66,Engineer,
      Employee67,Engineer,
      Employee68,Engineer,
      Employee69,Engineer,
      Employee70,Engineer,
      Employee71,Engineer,
      Employee72,Engineer,
      Employee73,Engineer,
      Employee74,Engineer,
      Employee75,Engineer,
      Employee76,Engineer,
      Employee77,Engineer,
      Employee78,Engineer,
      Employee79,Engineer,
      Employee80,Engineer,
      Employee81,Engineer,
      Employee82,Engineer,
      Employee83,Engineer,
      Employee84,Engineer,
      Employee85,Engineer,
      Employee86,Engineer,
      Employee87,Engineer,
      Employee88,Engineer,
      Employee89,Engineer,
      Employee90,Engineer,
      Employee91,Engineer,
      Employee92,Engineer,
      Employee93,Engineer,
      Employee94,Engineer,
      Employee95,Engineer,
      Employee96,Engineer,
      Employee97,Engineer,
      Employee98,Engineer,
      Employee99,Engineer,
      Employee100,Engineer
    ]
  ]
)--- 