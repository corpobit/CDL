---users:[name|n:age|b:active|t:date:joined:Alice,30,true,2025-05-19,Bob,25,false,2025-05-20,Charlie,28,true,2025-05-18]---
