---cities:[name|t:geo:coords|n:pop:NewYork,[40.7128,-74.0060],8398748,Tokyo,[35.6762,139.6503],37400068]---
