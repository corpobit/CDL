---data:[name|n:age|"home address":Alice,30,"123 Main St, NY",Bob,,null,"first name"|"n:last number":Charlie,42]---
